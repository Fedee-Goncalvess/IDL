library verilog;
use verilog.vl_types.all;
entity decodificador_salida_vlg_vec_tst is
end decodificador_salida_vlg_vec_tst;
