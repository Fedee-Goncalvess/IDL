library verilog;
use verilog.vl_types.all;
entity comparador_12bits_vlg_vec_tst is
end comparador_12bits_vlg_vec_tst;
