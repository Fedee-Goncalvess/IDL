library verilog;
use verilog.vl_types.all;
entity comparador_1bit_vlg_vec_tst is
end comparador_1bit_vlg_vec_tst;
