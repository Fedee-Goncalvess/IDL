library verilog;
use verilog.vl_types.all;
entity UC_estados_vlg_sample_tst is
    port(
        Q0              : in     vl_logic;
        Q1              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end UC_estados_vlg_sample_tst;
