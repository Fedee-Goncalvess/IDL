library verilog;
use verilog.vl_types.all;
entity unidad_control_vlg_vec_tst is
end unidad_control_vlg_vec_tst;
