library verilog;
use verilog.vl_types.all;
entity UC_de_UC_vlg_vec_tst is
end UC_de_UC_vlg_vec_tst;
