library verilog;
use verilog.vl_types.all;
entity UC_de_UA_vlg_vec_tst is
end UC_de_UA_vlg_vec_tst;
