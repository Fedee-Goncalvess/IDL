library verilog;
use verilog.vl_types.all;
entity UC_detector_fin_vlg_vec_tst is
end UC_detector_fin_vlg_vec_tst;
