library verilog;
use verilog.vl_types.all;
entity UC_detector_fin_vlg_check_tst is
    port(
        FIN             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end UC_detector_fin_vlg_check_tst;
