library verilog;
use verilog.vl_types.all;
entity conversorCA2_vlg_vec_tst is
end conversorCA2_vlg_vec_tst;
