library verilog;
use verilog.vl_types.all;
entity sumador_12bits_serie_vlg_vec_tst is
end sumador_12bits_serie_vlg_vec_tst;
