library verilog;
use verilog.vl_types.all;
entity UC_estados_vlg_vec_tst is
end UC_estados_vlg_vec_tst;
