library verilog;
use verilog.vl_types.all;
entity circuito_principal_bloque_vlg_vec_tst is
end circuito_principal_bloque_vlg_vec_tst;
